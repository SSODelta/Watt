module mux_2to1(Y, A, B, sel);
assign or__17__n_sel = (_17_ | (~ sel));
assign or__11__n_A0'h0 = (_11_ | (~ A[0]));
assign or__12__n_B0'h0 = (_12_ | (~ B[0]));
assign or__13__n_A1'h1 = (_13_ | (~ A[1]));
assign or__14__n_B1'h1 = (_14_ | (~ B[1]));
assign or__15__n__2_1'h1 = (_15_ | (~ _2_[1]));
assign or__16__n__1_0'h0 = (_16_ | (~ _1_[0]));
assign or__09__and_sel__0_1'h1 = (_09_ | (sel & _0_[1]));
assign or__10__and__17___2_1'h1 = (_10_ | (_17_ & _2_[1]));
assign or_Y1'h1_or__09___10_ = (Y[1] | (_09_ | _10_));
assign or__03__and__11__B0'h0 = (_03_ | (_11_ & B[0]));
assign or__04__and_A0'h0__12_ = (_04_ | (A[0] & _12_));
assign or_Y0'h0_or__03___04_ = (Y[0] | (_03_ | _04_));
assign or__05__and__13__B1'h1 = (_05_ | (_13_ & B[1]));
assign or__06__and_A1'h1__14_ = (_06_ | (A[1] & _14_));
assign or__2_1'h1_or__05___06_ = (_2_[1] | (_05_ | _06_));
assign or__07__and__15___1_0'h0 = (_07_ | (_15_ & _1_[0]));
assign or__08__and__2_1'h1__16_ = (_08_ | (_2_[1] & _16_));
assign or__0_1'h1_or__07___08_ = (_0_[1] | (_07_ | _08_));
assign or__1_0'h0_and_A0'h0_B0'h0 = (_1_[0] | (A[0] & B[0]));
endmodule
